module mux8tb;
reg i1,i2,i3,i4,i5,i6,i7,i8;
reg [2:0]s;
wire y;
mux8 dut(i1,i2,i3,i4,i5,i6,i7,i8,s,y);
initial begin
s=3'b000;i1=0;i2=0;i3=0;i4=0;i5=0;i6=0;i7=0;i8=0;
#10 i1=1;
#10 s=3'b001;i1=0;i2=0;i3=0;i4=0;i5=0;i6=0;i7=0;i8=0;
#10 i2=1;
#10 s=3'b010;i1=0;i2=0;i3=0;i4=0;i5=0;i6=0;i7=0;i8=0;
#10 i3=1;
#10 s=3'b011;i1=0;i2=0;i3=0;i4=0;i5=0;i6=0;i7=0;i8=0;
#10 i4=1;
#10 s=3'b100;i1=0;i2=0;i3=0;i4=0;i5=0;i6=0;i7=0;i8=0;
#10 i5=1;
#10 s=3'b101;i1=0;i2=0;i3=0;i4=0;i5=0;i6=0;i7=0;i8=0;
#10 i6=1;
#10 s=3'b110;i1=0;i2=0;i3=0;i4=0;i5=0;i6=0;i7=0;i8=0;
#10 i7=1;
#10 s=3'b111;i1=0;i2=0;i3=0;i4=0;i5=0;i6=0;i7=0;i8=0;
#10 i8=1;
#10 $finish();
end
endmodule